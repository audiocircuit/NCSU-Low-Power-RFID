library verilog;
use verilog.vl_types.all;
entity testbench1 is
end testbench1;
