module decode(
  input 




  );
