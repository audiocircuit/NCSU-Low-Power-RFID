library verilog;
use verilog.vl_types.all;
entity testbech is
end testbech;
