library verilog;
use verilog.vl_types.all;
entity tri_state_buffer_testbench is
end tri_state_buffer_testbench;
