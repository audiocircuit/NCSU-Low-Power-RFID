library verilog;
use verilog.vl_types.all;
entity I2C_testbench is
end I2C_testbench;
